module test
endmodule